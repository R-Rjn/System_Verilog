module prg(output bit [7:0] value);
  initial begin
    value<=20;
  end
endmodule
